module Tutorial(
);

// Welcome to Arctic Fox! In the first step, we will describe the code structure of an Automation. 
// It was important to us that Automations could be compiled by typical industry standard tools. 
// Therefore, to enable Automations to live within Verilog, we created them to be contained within
// comments. The following would be an Automation named ShiftReg, except that there would not be 
// a space between the * and either the [ or ]. 

/* [ShiftReg] */

// 1) Create an Automation with the name ShiftReg below. Do it  by typing the line above without a
//    space between the * and [ or ].


// If done correctly, it should look like the line below. The [ and ] should be grey, the /* and */
// should not be seen, and the ShiftReg should be bold. As the following: 
/*[ShiftReg]*/

// We got tired of having to type the Automation syntax constantly, so we made a shortcut. Start the 
// next tutorial to learn how to insert Automations easier.  

// To move between tutorials, you need to commit and changes and checkout the next tutorial step. For
// example, you need to add all 

endmodule